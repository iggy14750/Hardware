ENTITY DispBin IS
    PORT(
            
    );
END DispBin;

